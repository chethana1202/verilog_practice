module decoder4_10(D,Y);

input [3:0] D;
output reg [9:0] Y;

always@(*)
begin
    case(D)
    4'b0000: Y = 10'b0000000001;
    4'b0001: Y = 10'b0000000010;
    4'b0010: Y = 10'b0000000100;
    4'b0011: Y = 10'b0000001000;
    4'b0100: Y = 10'b0000010000;
    4'b0101: Y = 10'b0000100000;
    4'b0110: Y = 10'b0001000000;
    4'b0111: Y = 10'b0010000000;
    4'b1000: Y = 10'b0100000000;
    4'b1001: Y = 10'b1000000000;
    default: Y = 10'b0000000000;
    endcase
end

endmodule
